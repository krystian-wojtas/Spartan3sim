`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date:    19:22:47 08/18/2013
// Design Name:
// Module Name:    Sync
// Project Name:
// Target Devices:
// Tool versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////

module Sync (
        input  CLK50MHZ,
        input  RST,
        // vga interface
        output VGA_HSYNC,
        output VGA_VSYNC,
        // tick for next pixel
        output [10:0] x,
        output [10:0] y,
        output displaying
);

	localparam [10:0] H_S  = 2*800;
	localparam [ 1:0] H_FP = 2*16;
	localparam [ 7:0] H_PW = 2*96;
	localparam [ 6:0] H_BP = 2*48;
	localparam [ 9:0] V_S  = 521;
	localparam [ 1:0] V_PW = 2;
	localparam [ 3:0] V_FP = 10;
	localparam [ 4:0] V_BP = 29;

        wire [10:0] i;
        wire        h;
        Counter #(
                .MAX(H_S)
        ) Counter_h (
                .CLKB(CLK50MHZ),
                // counter
                .en(1'b1),
                .rst(RST),
                .sig(1'b1), // count all CLK50MHZ ticks
                .cnt(i),
                .full(h)
        );

        wire [9:0] j;
        Counter #(
                .MAX(V_S)
        ) Counter_v (
                .CLKB(CLK50MHZ),
                // counter
                .en(1'b1),
                .rst(RST),
                .sig(h), // count h sync
                .cnt(j)
        );

        assign displaying = (
            i >= H_PW + H_BP &&
            i <  H_S  - H_FP &&
            j >= V_BP + V_FP &&
            j <  V_S  - V_PW
        );

        assign VGA_HSYNC = (i > 96);
        assign VGA_VSYNC = (j > 2);

        assign x = i - 144;
        assign y = j - 39;

endmodule
